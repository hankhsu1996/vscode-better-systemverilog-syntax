// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.10--celldefine-basic-1
:description: Test
:tags: 22.10
:type: preprocessing
*/
`celldefine
//<----------- keyword.control.celldefine.sv
`endcelldefine
//<------------- keyword.control.endcelldefine.sv
