// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'property' token, color it immediately.

property
//<------- storage.type.property.sv
