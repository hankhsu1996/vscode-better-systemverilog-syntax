// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'interface' token, color it immediately.

interface
//<------ storage.type.interface.sv
