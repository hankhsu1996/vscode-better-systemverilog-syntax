// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: event
:description: event type tests
:tags: 6.17
*/
module top();
  event a;
//^^^^^ entity.name.type.event.sv
endmodule
