// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'macromodule' token, color it immediately.

macromodule
//<----------- storage.type.macromodule.sv
