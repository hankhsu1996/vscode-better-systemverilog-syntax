// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.11--pragma-invalid
:description: Test
:should_fail_because: The pragma specification is identified by the pragma_name, which follows the `pragma directive.
:tags: 22.11
:type: preprocessing
*/
`pragma
//<------- keyword.control.pragma.sv
