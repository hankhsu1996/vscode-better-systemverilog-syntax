// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'class' token, color it immediately.

class
//<------ storage.type.class.sv
