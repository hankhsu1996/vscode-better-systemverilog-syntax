// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'config' token, color it immediately.

config
//<------- storage.type.config.sv
