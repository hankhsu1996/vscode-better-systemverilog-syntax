// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'task' token, color it immediately.

task
//<------- storage.type.task.sv
