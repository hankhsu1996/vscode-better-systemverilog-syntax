// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'function' token, color it immediately.

function
//<------- storage.type.function.sv
