// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: chandle
:description: chandle type tests
:tags: 6.14
*/
module top();
  chandle a;
//^^^^^^^ entity.name.type.chandle.sv
endmodule
