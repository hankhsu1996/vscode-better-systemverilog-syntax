// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'module' token, color it immediately.

module
//<------ storage.type.module.sv
