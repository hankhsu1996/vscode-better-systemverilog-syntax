// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: array_addressing_sim
:description: array addressing simulation test
:type: simulation elaboration parsing
:tags: 11.5.2
*/
module top();
logic [7:0] mem [0:1023];
logic [7:0] a;

initial begin
  mem[123] = 125;
//   ^^^^^ meta.dimension.sv
//    ^^^ constant.numeric.integer.sv
  a = mem[123];
//       ^^^^^ meta.dimension.sv
//        ^^^ constant.numeric.integer.sv
  $display(":assert: (125 == %d)", a);
end

endmodule
