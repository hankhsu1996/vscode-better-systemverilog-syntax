// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: basic-unpacked
:description: Test unpacked arrays support
:tags: 7.4.2 7.4
*/
module top ();

bit _bit [7:0];
logic _logic [7:0];
reg _reg [7:0];

endmodule
