// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: manually_seeding_randomize_0
:description: manually seeding randomize test
:tags: 18.15
*/

class a;
    rand int x;
    function new (int seed);
        this.srandom(seed);
//           ^^^^^^^ entity.name.function.sv
    endfunction
endclass
