// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: nettype
:description: user-defined nettype tests
:tags: 6.6.7
*/
module top();
  nettype real real_net;
//^^^^^^^ keyword.control.nettype.sv
//        ^^^^ entity.name.type.sv
//             ^^^^^^^^ entity.name.type.sv
endmodule
