// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.9--unconnected_drive-basic-2
:description: Test
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull1
//<------------------ keyword.control.unconnected-drive.sv
//                 ^^^^^ storage.modifier.pull1.sv
