// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'interface class' token, color it immediately.

interface class
//<--------- storage.type.interface.sv
//        ^^^^^ storage.type.class.sv
