// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'sequence' token, color it immediately.

sequence
//<------- storage.type.sequence.sv
