// SYNTAX TEST "source-text.sv"

module Test;

<<<<<<< HEAD
  adder a1(
//^^^^^ entity.name.type.sv
//      ^^ variable.other.sv
    .a(a),
    .b(b)
  );
=======
  adder a2(
//^^^^^ entity.name.type.sv
//      ^^ variable.other.sv
    .a(a),
    .b(b)
  );
>>>>>>> branch-a
endmodule
