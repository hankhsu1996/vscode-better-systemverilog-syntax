// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.5.1--define_expansion_22
:description: Test
:tags: 22.5.1
:type: preprocessing
*/
`define max(a,b)((a) > (b) ? (a) : (b))
//                ^ variable.other.sv
//                   ^ keyword.operator.binary.sv
//                      ^ variable.other.sv
//                         ^ keyword.operator.ternary.sv
//                            ^ variable.other.sv
//                               ^ punctuation.separator.colon.sv
//                                  ^ variable.other.sv
