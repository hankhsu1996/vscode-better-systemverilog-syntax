// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.12--line-illegal-5
:description: Missing filename
:should_fail_because: Missing filename
:tags: 22.12
:type: preprocessing
*/
`line 1
//<----- keyword.control.line.sv
//    ^ constant.numeric.integer.sv
