// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'program' token, color it immediately.

program
//<------ storage.type.program.sv
