// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: 22.8--default_nettype
:description: Test
:tags: 22.8
:type: preprocessing
*/
`default_nettype wire
//<---------------- keyword.control.default-nettype.sv
//               ^^^^ entity.name.type.wire.sv
