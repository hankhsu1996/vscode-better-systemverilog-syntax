// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'covergroup' token, color it immediately.

covergroup
//<---------- storage.type.covergroup.sv
