// SYNTAX TEST "source-text.sv"
//
// Original source code by The SymbiFlow Authors under ISC License.
// Modifications by Shou-Li Hsu under MIT License.
// For full license information, see LICENSE file in the project root.
//
// vscode-tmgrammar-test annotations added by Shou-Li Hsu


/*
:name: string
:description: string type tests
:tags: 6.16
*/
module top();
  string a;
//^^^^^^ entity.name.type.string.sv
endmodule
