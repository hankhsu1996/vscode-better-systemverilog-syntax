// SYNTAX TEST "source-text.sv"

// Fail safe test: when we only have the 'package' token, color it immediately.

package
//<------- storage.type.package.sv
